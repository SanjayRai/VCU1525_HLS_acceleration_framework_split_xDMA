// Sanjay Rai (sanjay.d.rai@gmail.com)
//
`timescale 1 ps / 1 ps

module role_NORTH (
  input AXI_RESET_N,
  input CLK_IN_125M,
  input CLK_IN_250,
  input CLK_IN_PROG,
  input c0_sys_clk_n,
  input c0_sys_clk_p,
  input c2_sys_clk_n,
  input c2_sys_clk_p,
  input c3_sys_clk_n,
  input c3_sys_clk_p,
  output c0_ddr4_act_n,
  output [16:0]c0_ddr4_adr,
  output [1:0]c0_ddr4_ba,
  output [1:0]c0_ddr4_bg,
  output [0:0]c0_ddr4_ck_c,
  output [0:0]c0_ddr4_ck_t,
  output [0:0]c0_ddr4_cke,
  output [0:0]c0_ddr4_cs_n,
  inout [71:0]c0_ddr4_dq,
  inout [17:0]c0_ddr4_dqs_c,
  inout [17:0]c0_ddr4_dqs_t,
  output [0:0]c0_ddr4_odt,
  output c0_ddr4_par,
  output c0_ddr4_reset_n,
  output c0_init_calib_complete,
  output c2_ddr4_act_n,
  output [16:0]c2_ddr4_adr,
  output [1:0]c2_ddr4_ba,
  output [1:0]c2_ddr4_bg,
  output [0:0]c2_ddr4_ck_c,
  output [0:0]c2_ddr4_ck_t,
  output [0:0]c2_ddr4_cke,
  output [0:0]c2_ddr4_cs_n,
  inout [71:0]c2_ddr4_dq,
  inout [17:0]c2_ddr4_dqs_c,
  inout [17:0]c2_ddr4_dqs_t,
  output [0:0]c2_ddr4_odt,
  output c2_ddr4_par,
  output c2_ddr4_reset_n,
  output c2_init_calib_complete,
  output c3_ddr4_act_n,
  output [16:0]c3_ddr4_adr,
  output [1:0]c3_ddr4_ba,
  output [1:0]c3_ddr4_bg,
  output [0:0]c3_ddr4_ck_c,
  output [0:0]c3_ddr4_ck_t,
  output [0:0]c3_ddr4_cke,
  output [0:0]c3_ddr4_cs_n,
  inout [71:0]c3_ddr4_dq,
  inout [17:0]c3_ddr4_dqs_c,
  inout [17:0]c3_ddr4_dqs_t,
  output [0:0]c3_ddr4_odt,
  output c3_ddr4_par,
  output c3_ddr4_reset_n,
  output c3_init_calib_complete,
  output [31:0]ker_count,
  output ker_count_ap_vld,
  input sys_rst_ddr_0,
  input sys_rst_ddr_2,
  input sys_rst_ddr_3,
  srai_accel_AXI_MM_intfc.master M_AXI_NORTH_TO_STATIC,
  srai_accel_AXI_MM_intfc.slave S_AXI_FROM_STATIC,
  srai_accel_AXI_LITE_intfc.slave S_AXI_LITE_FROM_STATIC,
  input wire  S_BSCAN_bscanid_en,
  input wire  S_BSCAN_capture,
  input wire  S_BSCAN_drck,
  input wire  S_BSCAN_reset,
  input wire  S_BSCAN_runtest,
  input wire  S_BSCAN_sel,
  input wire  S_BSCAN_shift,
  input wire  S_BSCAN_tck,
  input wire  S_BSCAN_tdi,
  output wire S_BSCAN_tdo,
  input wire  S_BSCAN_tms,
  input wire  S_BSCAN_update
  );

  reg start_ker_r = 1'b0;
  reg start_ker_vld_r = 1'b0;


  HLS_PR_SDX_SRAI HLS_PR_0_i_NORTH
       (.AXI_RESET_N(AXI_RESET_N),
        .C0_SYS_CLK_clk_n(c0_sys_clk_n),
        .C0_SYS_CLK_clk_p(c0_sys_clk_p),
        .C2_SYS_CLK_clk_n(c2_sys_clk_n),
        .C2_SYS_CLK_clk_p(c2_sys_clk_p),
        .C3_SYS_CLK_clk_n(c3_sys_clk_n),
        .C3_SYS_CLK_clk_p(c3_sys_clk_p),
        .CLK_IN_125M(CLK_IN_125M),
        .CLK_IN_250(CLK_IN_250),
        .CLK_IN_PROG(CLK_IN_PROG),
        .M_AXI_TO_STATIC_araddr(M_AXI_NORTH_TO_STATIC.AXI_araddr),
        .M_AXI_TO_STATIC_arburst(M_AXI_NORTH_TO_STATIC.AXI_arburst),
        .M_AXI_TO_STATIC_arcache(M_AXI_NORTH_TO_STATIC.AXI_arcache),
        .M_AXI_TO_STATIC_arid(M_AXI_NORTH_TO_STATIC.AXI_arid[4:0]),
        .M_AXI_TO_STATIC_arlen(M_AXI_NORTH_TO_STATIC.AXI_arlen),
        .M_AXI_TO_STATIC_arlock(M_AXI_NORTH_TO_STATIC.AXI_arlock),
        .M_AXI_TO_STATIC_arprot(M_AXI_NORTH_TO_STATIC.AXI_arprot),
        .M_AXI_TO_STATIC_arqos(M_AXI_NORTH_TO_STATIC.AXI_arqos),
        .M_AXI_TO_STATIC_arready(M_AXI_NORTH_TO_STATIC.AXI_arready),
        .M_AXI_TO_STATIC_arregion(M_AXI_NORTH_TO_STATIC.AXI_arregion),
        .M_AXI_TO_STATIC_arsize(M_AXI_NORTH_TO_STATIC.AXI_arsize),
        .M_AXI_TO_STATIC_arvalid(M_AXI_NORTH_TO_STATIC.AXI_arvalid),
        .M_AXI_TO_STATIC_awaddr(M_AXI_NORTH_TO_STATIC.AXI_awaddr),
        .M_AXI_TO_STATIC_awburst(M_AXI_NORTH_TO_STATIC.AXI_awburst),
        .M_AXI_TO_STATIC_awcache(M_AXI_NORTH_TO_STATIC.AXI_awcache),
        .M_AXI_TO_STATIC_awid(M_AXI_NORTH_TO_STATIC.AXI_awid[4:0]),
        .M_AXI_TO_STATIC_awlen(M_AXI_NORTH_TO_STATIC.AXI_awlen),
        .M_AXI_TO_STATIC_awlock(M_AXI_NORTH_TO_STATIC.AXI_awlock),
        .M_AXI_TO_STATIC_awprot(M_AXI_NORTH_TO_STATIC.AXI_awprot),
        .M_AXI_TO_STATIC_awqos(M_AXI_NORTH_TO_STATIC.AXI_awqos),
        .M_AXI_TO_STATIC_awready(M_AXI_NORTH_TO_STATIC.AXI_awready),
        .M_AXI_TO_STATIC_awregion(M_AXI_NORTH_TO_STATIC.AXI_awregion),
        .M_AXI_TO_STATIC_awsize(M_AXI_NORTH_TO_STATIC.AXI_awsize),
        .M_AXI_TO_STATIC_awvalid(M_AXI_NORTH_TO_STATIC.AXI_awvalid),
        .M_AXI_TO_STATIC_bid(M_AXI_NORTH_TO_STATIC.AXI_bid[4:0]),
        .M_AXI_TO_STATIC_bready(M_AXI_NORTH_TO_STATIC.AXI_bready),
        .M_AXI_TO_STATIC_bresp(M_AXI_NORTH_TO_STATIC.AXI_bresp),
        .M_AXI_TO_STATIC_bvalid(M_AXI_NORTH_TO_STATIC.AXI_bvalid),
        .M_AXI_TO_STATIC_rdata(M_AXI_NORTH_TO_STATIC.AXI_rdata),
        .M_AXI_TO_STATIC_rid(M_AXI_NORTH_TO_STATIC.AXI_rid[4:0]),
        .M_AXI_TO_STATIC_rlast(M_AXI_NORTH_TO_STATIC.AXI_rlast),
        .M_AXI_TO_STATIC_rready(M_AXI_NORTH_TO_STATIC.AXI_rready),
        .M_AXI_TO_STATIC_rresp(M_AXI_NORTH_TO_STATIC.AXI_rresp),
        .M_AXI_TO_STATIC_rvalid(M_AXI_NORTH_TO_STATIC.AXI_rvalid),
        .M_AXI_TO_STATIC_wdata(M_AXI_NORTH_TO_STATIC.AXI_wdata),
        .M_AXI_TO_STATIC_wlast(M_AXI_NORTH_TO_STATIC.AXI_wlast),
        .M_AXI_TO_STATIC_wready(M_AXI_NORTH_TO_STATIC.AXI_wready),
        .M_AXI_TO_STATIC_wstrb(M_AXI_NORTH_TO_STATIC.AXI_wstrb),
        .M_AXI_TO_STATIC_wvalid(M_AXI_NORTH_TO_STATIC.AXI_wvalid),
        .S_AXI_FROM_STATIC_araddr(S_AXI_FROM_STATIC.AXI_araddr),
        .S_AXI_FROM_STATIC_arburst(S_AXI_FROM_STATIC.AXI_arburst),
        .S_AXI_FROM_STATIC_arcache(S_AXI_FROM_STATIC.AXI_arcache),
        .S_AXI_FROM_STATIC_arid(S_AXI_FROM_STATIC.AXI_arid[3:0]),
        .S_AXI_FROM_STATIC_arlen(S_AXI_FROM_STATIC.AXI_arlen),
        .S_AXI_FROM_STATIC_arlock(S_AXI_FROM_STATIC.AXI_arlock),
        .S_AXI_FROM_STATIC_arprot(S_AXI_FROM_STATIC.AXI_arprot),
        .S_AXI_FROM_STATIC_arqos(S_AXI_FROM_STATIC.AXI_arqos),
        .S_AXI_FROM_STATIC_arready(S_AXI_FROM_STATIC.AXI_arready),
        .S_AXI_FROM_STATIC_arregion(S_AXI_FROM_STATIC.AXI_arregion),
        .S_AXI_FROM_STATIC_arsize(S_AXI_FROM_STATIC.AXI_arsize),
        .S_AXI_FROM_STATIC_arvalid(S_AXI_FROM_STATIC.AXI_arvalid),
        .S_AXI_FROM_STATIC_awaddr(S_AXI_FROM_STATIC.AXI_awaddr),
        .S_AXI_FROM_STATIC_awburst(S_AXI_FROM_STATIC.AXI_awburst),
        .S_AXI_FROM_STATIC_awcache(S_AXI_FROM_STATIC.AXI_awcache),
        .S_AXI_FROM_STATIC_awid(S_AXI_FROM_STATIC.AXI_awid[3:0]),
        .S_AXI_FROM_STATIC_awlen(S_AXI_FROM_STATIC.AXI_awlen),
        .S_AXI_FROM_STATIC_awlock(S_AXI_FROM_STATIC.AXI_awlock),
        .S_AXI_FROM_STATIC_awprot(S_AXI_FROM_STATIC.AXI_awprot),
        .S_AXI_FROM_STATIC_awqos(S_AXI_FROM_STATIC.AXI_awqos),
        .S_AXI_FROM_STATIC_awready(S_AXI_FROM_STATIC.AXI_awready),
        .S_AXI_FROM_STATIC_awregion(S_AXI_FROM_STATIC.AXI_awregion),
        .S_AXI_FROM_STATIC_awsize(S_AXI_FROM_STATIC.AXI_awsize),
        .S_AXI_FROM_STATIC_awvalid(S_AXI_FROM_STATIC.AXI_awvalid),
        .S_AXI_FROM_STATIC_bid(S_AXI_FROM_STATIC.AXI_bid[3:0]),
        .S_AXI_FROM_STATIC_bready(S_AXI_FROM_STATIC.AXI_bready),
        .S_AXI_FROM_STATIC_bresp(S_AXI_FROM_STATIC.AXI_bresp),
        .S_AXI_FROM_STATIC_bvalid(S_AXI_FROM_STATIC.AXI_bvalid),
        .S_AXI_FROM_STATIC_rdata(S_AXI_FROM_STATIC.AXI_rdata),
        .S_AXI_FROM_STATIC_rid(S_AXI_FROM_STATIC.AXI_rid[3:0]),
        .S_AXI_FROM_STATIC_rlast(S_AXI_FROM_STATIC.AXI_rlast),
        .S_AXI_FROM_STATIC_rready(S_AXI_FROM_STATIC.AXI_rready),
        .S_AXI_FROM_STATIC_rresp(S_AXI_FROM_STATIC.AXI_rresp),
        .S_AXI_FROM_STATIC_rvalid(S_AXI_FROM_STATIC.AXI_rvalid),
        .S_AXI_FROM_STATIC_wdata(S_AXI_FROM_STATIC.AXI_wdata),
        .S_AXI_FROM_STATIC_wlast(S_AXI_FROM_STATIC.AXI_wlast),
        .S_AXI_FROM_STATIC_wready(S_AXI_FROM_STATIC.AXI_wready),
        .S_AXI_FROM_STATIC_wstrb(S_AXI_FROM_STATIC.AXI_wstrb),
        .S_AXI_FROM_STATIC_wvalid(S_AXI_FROM_STATIC.AXI_wvalid),
        .S_AXI_LITE_FROM_STATIC_araddr(S_AXI_LITE_FROM_STATIC.AXI_LITE_araddr),
        .S_AXI_LITE_FROM_STATIC_arprot(S_AXI_LITE_FROM_STATIC.AXI_LITE_arprot),
        .S_AXI_LITE_FROM_STATIC_arready(S_AXI_LITE_FROM_STATIC.AXI_LITE_arready),
        .S_AXI_LITE_FROM_STATIC_arvalid(S_AXI_LITE_FROM_STATIC.AXI_LITE_arvalid),
        .S_AXI_LITE_FROM_STATIC_awaddr(S_AXI_LITE_FROM_STATIC.AXI_LITE_awaddr),
        .S_AXI_LITE_FROM_STATIC_awprot(S_AXI_LITE_FROM_STATIC.AXI_LITE_awprot),
        .S_AXI_LITE_FROM_STATIC_awready(S_AXI_LITE_FROM_STATIC.AXI_LITE_awready),
        .S_AXI_LITE_FROM_STATIC_awvalid(S_AXI_LITE_FROM_STATIC.AXI_LITE_awvalid),
        .S_AXI_LITE_FROM_STATIC_bready(S_AXI_LITE_FROM_STATIC.AXI_LITE_bready),
        .S_AXI_LITE_FROM_STATIC_bresp(S_AXI_LITE_FROM_STATIC.AXI_LITE_bresp),
        .S_AXI_LITE_FROM_STATIC_bvalid(S_AXI_LITE_FROM_STATIC.AXI_LITE_bvalid),
        .S_AXI_LITE_FROM_STATIC_rdata(S_AXI_LITE_FROM_STATIC.AXI_LITE_rdata),
        .S_AXI_LITE_FROM_STATIC_rready(S_AXI_LITE_FROM_STATIC.AXI_LITE_rready),
        .S_AXI_LITE_FROM_STATIC_rresp(S_AXI_LITE_FROM_STATIC.AXI_LITE_rresp),
        .S_AXI_LITE_FROM_STATIC_rvalid(S_AXI_LITE_FROM_STATIC.AXI_LITE_rvalid),
        .S_AXI_LITE_FROM_STATIC_wdata(S_AXI_LITE_FROM_STATIC.AXI_LITE_wdata),
        .S_AXI_LITE_FROM_STATIC_wready(S_AXI_LITE_FROM_STATIC.AXI_LITE_wready),
        .S_AXI_LITE_FROM_STATIC_wstrb(S_AXI_LITE_FROM_STATIC.AXI_LITE_wstrb),
        .S_AXI_LITE_FROM_STATIC_wvalid(S_AXI_LITE_FROM_STATIC.AXI_LITE_wvalid),
        .c0_ddr4_act_n(c0_ddr4_act_n),
        .c0_ddr4_adr(c0_ddr4_adr),
        .c0_ddr4_ba(c0_ddr4_ba),
        .c0_ddr4_bg(c0_ddr4_bg),
        .c0_ddr4_ck_c(c0_ddr4_ck_c),
        .c0_ddr4_ck_t(c0_ddr4_ck_t),
        .c0_ddr4_cke(c0_ddr4_cke),
        .c0_ddr4_cs_n(c0_ddr4_cs_n),
        .c0_ddr4_dq(c0_ddr4_dq),
        .c0_ddr4_dqs_c(c0_ddr4_dqs_c),
        .c0_ddr4_dqs_t(c0_ddr4_dqs_t),
        .c0_ddr4_odt(c0_ddr4_odt),
        .c0_ddr4_par(c0_ddr4_par),
        .c0_ddr4_reset_n(c0_ddr4_reset_n),
        .c0_init_calib_complete(c0_init_calib_complete),
        .c2_ddr4_act_n(c2_ddr4_act_n),
        .c2_ddr4_adr(c2_ddr4_adr),
        .c2_ddr4_ba(c2_ddr4_ba),
        .c2_ddr4_bg(c2_ddr4_bg),
        .c2_ddr4_ck_c(c2_ddr4_ck_c),
        .c2_ddr4_ck_t(c2_ddr4_ck_t),
        .c2_ddr4_cke(c2_ddr4_cke),
        .c2_ddr4_cs_n(c2_ddr4_cs_n),
        .c2_ddr4_dq(c2_ddr4_dq),
        .c2_ddr4_dqs_c(c2_ddr4_dqs_c),
        .c2_ddr4_dqs_t(c2_ddr4_dqs_t),
        .c2_ddr4_odt(c2_ddr4_odt),
        .c2_ddr4_par(c2_ddr4_par),
        .c2_ddr4_reset_n(c2_ddr4_reset_n),
        .c2_init_calib_complete(c2_init_calib_complete),
        .c3_ddr4_act_n(c3_ddr4_act_n),
        .c3_ddr4_adr(c3_ddr4_adr),
        .c3_ddr4_ba(c3_ddr4_ba),
        .c3_ddr4_bg(c3_ddr4_bg),
        .c3_ddr4_ck_c(c3_ddr4_ck_c),
        .c3_ddr4_ck_t(c3_ddr4_ck_t),
        .c3_ddr4_cke(c3_ddr4_cke),
        .c3_ddr4_cs_n(c3_ddr4_cs_n),
        .c3_ddr4_dq(c3_ddr4_dq),
        .c3_ddr4_dqs_c(c3_ddr4_dqs_c),
        .c3_ddr4_dqs_t(c3_ddr4_dqs_t),
        .c3_ddr4_odt(c3_ddr4_odt),
        .c3_ddr4_par(c3_ddr4_par),
        .c3_ddr4_reset_n(c3_ddr4_reset_n),
        .c3_init_calib_complete(c3_init_calib_complete),
        .ker_count(ker_count),
        .ker_count_ap_vld(ker_count_ap_vld),
        .sys_rst_ddr_0(sys_rst_ddr_0),
        .sys_rst_ddr_2(sys_rst_ddr_2),
        .sys_rst_ddr_3(sys_rst_ddr_3));

//ila_0 U_ila_0 (
//	.clk(CLK_IN_PROG), // input wire clk
//	.probe0({start_ker_vld_r, start_ker_r}) // input wire [0:0] probe0
//);

debug_bridge_PR U_debug_bridge_PR (
  .clk(CLK_IN_125M),                                // input wire clk
  .S_BSCAN_bscanid_en(S_BSCAN_bscanid_en),  // input wire s_bscan_bscanid_en
  .S_BSCAN_capture(S_BSCAN_capture),        // input wire s_bscan_capture
  .S_BSCAN_drck(S_BSCAN_drck),              // input wire s_bscan_drck
  .S_BSCAN_reset(S_BSCAN_reset),            // input wire s_bscan_reset
  .S_BSCAN_runtest(S_BSCAN_runtest),        // input wire s_bscan_runtest
  .S_BSCAN_sel(S_BSCAN_sel),                // input wire s_bscan_sel
  .S_BSCAN_shift(S_BSCAN_shift),            // input wire s_bscan_shift
  .S_BSCAN_tck(S_BSCAN_tck),                // input wire s_bscan_tck
  .S_BSCAN_tdi(S_BSCAN_tdi),                // input wire s_bscan_tdi
  .S_BSCAN_tdo(S_BSCAN_tdo),                // output wire s_bscan_tdo
  .S_BSCAN_tms(S_BSCAN_tms),                // input wire s_bscan_tms
  .S_BSCAN_update(S_BSCAN_update)          // input wire s_bscan_update
);

endmodule
