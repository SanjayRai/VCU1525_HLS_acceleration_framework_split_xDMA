// Sanjay Rai (sanjay.d.rai@gmail.com)
//
`timescale 1 ps / 1 ps

module VU9P_AXI_ICAP_PR_DESIGN_top (
  input c0_sys_clk_n,
  input c0_sys_clk_p,
  input c1_sys_clk_n,
  input c1_sys_clk_p,
  input c2_sys_clk_n,
  input c2_sys_clk_p,
  input c3_sys_clk_n,
  input c3_sys_clk_p,

  output c0_ddr4_act_n,
  output [16:0]c0_ddr4_adr,
  output [1:0]c0_ddr4_ba,
  output [1:0]c0_ddr4_bg,
  output [0:0]c0_ddr4_ck_c,
  output [0:0]c0_ddr4_ck_t,
  output [0:0]c0_ddr4_cke,
  output [0:0]c0_ddr4_cs_n,
  inout [71:0]c0_ddr4_dq,
  inout [17:0]c0_ddr4_dqs_c,
  inout [17:0]c0_ddr4_dqs_t,
  output [0:0]c0_ddr4_odt,
  output c0_ddr4_par,
  output c0_ddr4_reset_n,

  output c1_ddr4_act_n,
  output [16:0]c1_ddr4_adr,
  output [1:0]c1_ddr4_ba,
  output [1:0]c1_ddr4_bg,
  output [0:0]c1_ddr4_ck_c,
  output [0:0]c1_ddr4_ck_t,
  output [0:0]c1_ddr4_cke,
  output [0:0]c1_ddr4_cs_n,
  inout [71:0]c1_ddr4_dq,
  inout [17:0]c1_ddr4_dqs_c,
  inout [17:0]c1_ddr4_dqs_t,
  output [0:0]c1_ddr4_odt,
  output c1_ddr4_par,
  output c1_ddr4_reset_n,
  output c2_ddr4_act_n,
  output [16:0]c2_ddr4_adr,
  output [1:0]c2_ddr4_ba,
  output [1:0]c2_ddr4_bg,
  output [0:0]c2_ddr4_ck_c,
  output [0:0]c2_ddr4_ck_t,
  output [0:0]c2_ddr4_cke,
  output [0:0]c2_ddr4_cs_n,
  inout [71:0]c2_ddr4_dq,
  inout [17:0]c2_ddr4_dqs_c,
  inout [17:0]c2_ddr4_dqs_t,
  output [0:0]c2_ddr4_odt,
  output c2_ddr4_par,
  output c2_ddr4_reset_n,
  output c3_ddr4_act_n,
  output [16:0]c3_ddr4_adr,
  output [1:0]c3_ddr4_ba,
  output [1:0]c3_ddr4_bg,
  output [0:0]c3_ddr4_ck_c,
  output [0:0]c3_ddr4_ck_t,
  output [0:0]c3_ddr4_cke,
  output [0:0]c3_ddr4_cs_n,
  inout [71:0]c3_ddr4_dq,
  inout [17:0]c3_ddr4_dqs_c,
  inout [17:0]c3_ddr4_dqs_t,
  output [0:0]c3_ddr4_odt,
  output c3_ddr4_par,
  output c3_ddr4_reset_n,
  input [15:0]pcie_mgt_rxn,
  input [15:0]pcie_mgt_rxp,
  output [15:0]pcie_mgt_txn,
  output [15:0]pcie_mgt_txp,
  input         sys_clk_p,
  input         sys_clk_n,
  input         sys_rst_n );

  wire sys_rst_n_c;
  wire sys_clk;
  wire sys_clk_gt;
  wire clk_out_125M;
  wire clk_out_250M;
  wire clk_out_PROG;
  wire axi_reset_n_out;
  wire [31:0]ker_count;
  wire ker_count_ap_vld;
  wire c0_init_calib_complete;
  wire c2_init_calib_complete;
  wire c3_init_calib_complete;

  IBUF   sys_reset_n_ibuf (.O(sys_rst_n_c), .I(sys_rst_n));
  IBUFDS_GTE4 refclk_ibuf (.O(sys_clk_gt), .ODIV2(sys_clk), .I(sys_clk_p), .CEB(1'b0), .IB(sys_clk_n));

  srai_accel_AXI_MM_intfc AXI_MM_FROM_HLS_PR ();
  srai_accel_AXI_MM_intfc AXI_MM_TO_HLS_PR ();
  srai_accel_AXI_LITE_intfc M_AXI_LITE_TO_HLS_PR();

  shell_top U_shell_top (
        .C1_SYS_CLK_clk_n(c1_sys_clk_n),
        .C1_SYS_CLK_clk_p(c1_sys_clk_p),
        .DDR4_sys_rst(1'b0),
        .M_AXI_LITE_TO_HLS_PR_NORTH(M_AXI_LITE_TO_HLS_PR.master),
        .S_AXI_MM_FROM_HLS_PR_NORTH(AXI_MM_FROM_HLS_PR.slave),
        .M_AXI_MM_TO_HLS_PR_NORTH(AXI_MM_TO_HLS_PR.master),
        .axi_reset_n_out(axi_reset_n_out),
        .c1_ddr4_act_n(c1_ddr4_act_n),
        .c1_ddr4_adr(c1_ddr4_adr),
        .c1_ddr4_ba(c1_ddr4_ba),
        .c1_ddr4_bg(c1_ddr4_bg),
        .c1_ddr4_ck_c(c1_ddr4_ck_c),
        .c1_ddr4_ck_t(c1_ddr4_ck_t),
        .c1_ddr4_cke(c1_ddr4_cke),
        .c1_ddr4_cs_n(c1_ddr4_cs_n),
        .c1_ddr4_par(c1_ddr4_par),
        .c1_ddr4_dq(c1_ddr4_dq),
        .c1_ddr4_dqs_c(c1_ddr4_dqs_c),
        .c1_ddr4_dqs_t(c1_ddr4_dqs_t),
        .c1_ddr4_odt(c1_ddr4_odt),
        .c1_ddr4_reset_n(c1_ddr4_reset_n),
        .clk_out_125M(clk_out_125M),
        .clk_out_250M(clk_out_250M),
        .clk_out_PROG(clk_out_PROG),
        .ker_count(ker_count),
        .ker_count_ap_vld(ker_count_ap_vld),
        .c0_init_calib_complete(c0_init_calib_complete),
        .c2_init_calib_complete(c2_init_calib_complete),
        .c3_init_calib_complete(c3_init_calib_complete),
        .pcie_mgt_rxn(pcie_mgt_rxn),
        .pcie_mgt_rxp(pcie_mgt_rxp),
        .pcie_mgt_txn(pcie_mgt_txn),
        .pcie_mgt_txp(pcie_mgt_txp),
        .sys_clk(sys_clk),
        .sys_clk_gt(sys_clk_gt),
        .sys_rst_n(sys_rst_n_c));


  role_NORTH U_role_NORTH (
        .AXI_RESET_N(axi_reset_n_out),
        .CLK_IN_250(clk_out_250M),
        .CLK_IN_125M(clk_out_125M),
        .CLK_IN_PROG(clk_out_PROG),
        .c0_sys_clk_n(c0_sys_clk_n),
        .c0_sys_clk_p(c0_sys_clk_p),
        .c2_sys_clk_n(c2_sys_clk_n),
        .c2_sys_clk_p(c2_sys_clk_p),
        .c3_sys_clk_n(c3_sys_clk_n),
        .c3_sys_clk_p(c3_sys_clk_p),
        .c0_ddr4_act_n(c0_ddr4_act_n),
        .c0_ddr4_adr(c0_ddr4_adr),
        .c0_ddr4_ba(c0_ddr4_ba),
        .c0_ddr4_bg(c0_ddr4_bg),
        .c0_ddr4_ck_c(c0_ddr4_ck_c),
        .c0_ddr4_ck_t(c0_ddr4_ck_t),
        .c0_ddr4_cke(c0_ddr4_cke),
        .c0_ddr4_cs_n(c0_ddr4_cs_n),
        .c0_ddr4_dq(c0_ddr4_dq),
        .c0_ddr4_dqs_c(c0_ddr4_dqs_c),
        .c0_ddr4_dqs_t(c0_ddr4_dqs_t),
        .c0_ddr4_odt(c0_ddr4_odt),
        .c0_ddr4_par(c0_ddr4_par),
        .c0_ddr4_reset_n(c0_ddr4_reset_n),
        .c0_init_calib_complete(c0_init_calib_complete),
        .c2_ddr4_act_n(c2_ddr4_act_n),
        .c2_ddr4_adr(c2_ddr4_adr),
        .c2_ddr4_ba(c2_ddr4_ba),
        .c2_ddr4_bg(c2_ddr4_bg),
        .c2_ddr4_ck_c(c2_ddr4_ck_c),
        .c2_ddr4_ck_t(c2_ddr4_ck_t),
        .c2_ddr4_cke(c2_ddr4_cke),
        .c2_ddr4_cs_n(c2_ddr4_cs_n),
        .c2_ddr4_dq(c2_ddr4_dq),
        .c2_ddr4_dqs_c(c2_ddr4_dqs_c),
        .c2_ddr4_dqs_t(c2_ddr4_dqs_t),
        .c2_ddr4_odt(c2_ddr4_odt),
        .c2_ddr4_par(c2_ddr4_par),
        .c2_ddr4_reset_n(c2_ddr4_reset_n),
        .c2_init_calib_complete(c2_init_calib_complete),
        .c3_ddr4_act_n(c3_ddr4_act_n),
        .c3_ddr4_adr(c3_ddr4_adr),
        .c3_ddr4_ba(c3_ddr4_ba),
        .c3_ddr4_bg(c3_ddr4_bg),
        .c3_ddr4_ck_c(c3_ddr4_ck_c),
        .c3_ddr4_ck_t(c3_ddr4_ck_t),
        .c3_ddr4_cke(c3_ddr4_cke),
        .c3_ddr4_cs_n(c3_ddr4_cs_n),
        .c3_ddr4_dq(c3_ddr4_dq),
        .c3_ddr4_dqs_c(c3_ddr4_dqs_c),
        .c3_ddr4_dqs_t(c3_ddr4_dqs_t),
        .c3_ddr4_odt(c3_ddr4_odt),
        .c3_ddr4_par(c3_ddr4_par),
        .c3_ddr4_reset_n(c3_ddr4_reset_n),
        .c3_init_calib_complete(c3_init_calib_complete),
        .ker_count(ker_count),
        .ker_count_ap_vld(ker_count_ap_vld),
        .sys_rst_ddr_0(1'b0),
        .sys_rst_ddr_2(1'b0),
        .sys_rst_ddr_3(1'b0),
        .M_AXI_NORTH_TO_STATIC(AXI_MM_FROM_HLS_PR.master),
        .S_AXI_FROM_STATIC (AXI_MM_TO_HLS_PR.slave),
        .S_AXI_LITE_FROM_STATIC(M_AXI_LITE_TO_HLS_PR.slave),
        .S_BSCAN_bscanid_en(),
        .S_BSCAN_capture(),
        .S_BSCAN_drck(),
        .S_BSCAN_reset(),
        .S_BSCAN_runtest(),
        .S_BSCAN_sel(),
        .S_BSCAN_shift(),
        .S_BSCAN_tck(),
        .S_BSCAN_tdi(),
        .S_BSCAN_tdo(),
        .S_BSCAN_tms(),
        .S_BSCAN_update()
        );

endmodule
